-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Sun Nov 30 11:56:14 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY div_freq IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		rst :  IN  STD_LOGIC;
		clkOUT :  OUT  STD_LOGIC
	);
END div_freq;

ARCHITECTURE bdf_type OF div_freq IS 

SIGNAL	clkOUT_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_50 <= '1';



PROCESS(clk,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_56 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_56 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_56 <= SYNTHESIZED_WIRE_0;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_51,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_53 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_53 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_51)) THEN
	SYNTHESIZED_WIRE_53 <= SYNTHESIZED_WIRE_2;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_48 <= NOT(SYNTHESIZED_WIRE_52);



PROCESS(SYNTHESIZED_WIRE_52,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_51 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_51 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_51 <= SYNTHESIZED_WIRE_4;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_4 <= NOT(SYNTHESIZED_WIRE_51);



SYNTHESIZED_WIRE_2 <= NOT(SYNTHESIZED_WIRE_53);




PROCESS(SYNTHESIZED_WIRE_53,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_54 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_54 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_53)) THEN
	SYNTHESIZED_WIRE_54 <= SYNTHESIZED_WIRE_6;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_6 <= NOT(SYNTHESIZED_WIRE_54);



PROCESS(SYNTHESIZED_WIRE_54,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_55 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_55 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_54)) THEN
	SYNTHESIZED_WIRE_55 <= SYNTHESIZED_WIRE_8;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_8 <= NOT(SYNTHESIZED_WIRE_55);



PROCESS(SYNTHESIZED_WIRE_55,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_57 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_57 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_55)) THEN
	SYNTHESIZED_WIRE_57 <= SYNTHESIZED_WIRE_10;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_0 <= NOT(SYNTHESIZED_WIRE_56);



SYNTHESIZED_WIRE_10 <= NOT(SYNTHESIZED_WIRE_57);



PROCESS(SYNTHESIZED_WIRE_57,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_58 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_58 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_57)) THEN
	SYNTHESIZED_WIRE_58 <= SYNTHESIZED_WIRE_12;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_12 <= NOT(SYNTHESIZED_WIRE_58);



PROCESS(SYNTHESIZED_WIRE_58,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_59 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_59 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_58)) THEN
	SYNTHESIZED_WIRE_59 <= SYNTHESIZED_WIRE_14;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_14 <= NOT(SYNTHESIZED_WIRE_59);



PROCESS(SYNTHESIZED_WIRE_59,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_60 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_60 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_59)) THEN
	SYNTHESIZED_WIRE_60 <= SYNTHESIZED_WIRE_16;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_16 <= NOT(SYNTHESIZED_WIRE_60);



PROCESS(SYNTHESIZED_WIRE_60,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_61 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_61 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_60)) THEN
	SYNTHESIZED_WIRE_61 <= SYNTHESIZED_WIRE_18;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_18 <= NOT(SYNTHESIZED_WIRE_61);



PROCESS(SYNTHESIZED_WIRE_61,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_62 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_62 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_61)) THEN
	SYNTHESIZED_WIRE_62 <= SYNTHESIZED_WIRE_20;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_56,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_67 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_67 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_56)) THEN
	SYNTHESIZED_WIRE_67 <= SYNTHESIZED_WIRE_22;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_20 <= NOT(SYNTHESIZED_WIRE_62);



PROCESS(SYNTHESIZED_WIRE_62,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_63 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_63 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_62)) THEN
	SYNTHESIZED_WIRE_63 <= SYNTHESIZED_WIRE_24;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_24 <= NOT(SYNTHESIZED_WIRE_63);



PROCESS(SYNTHESIZED_WIRE_63,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_64 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_64 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_63)) THEN
	SYNTHESIZED_WIRE_64 <= SYNTHESIZED_WIRE_26;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_26 <= NOT(SYNTHESIZED_WIRE_64);



PROCESS(SYNTHESIZED_WIRE_64,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_65 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_65 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_64)) THEN
	SYNTHESIZED_WIRE_65 <= SYNTHESIZED_WIRE_28;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_28 <= NOT(SYNTHESIZED_WIRE_65);



PROCESS(SYNTHESIZED_WIRE_65,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_66 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_66 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_65)) THEN
	SYNTHESIZED_WIRE_66 <= SYNTHESIZED_WIRE_30;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_30 <= NOT(SYNTHESIZED_WIRE_66);



PROCESS(SYNTHESIZED_WIRE_66,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_68 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_68 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_66)) THEN
	SYNTHESIZED_WIRE_68 <= SYNTHESIZED_WIRE_32;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_22 <= NOT(SYNTHESIZED_WIRE_67);



SYNTHESIZED_WIRE_32 <= NOT(SYNTHESIZED_WIRE_68);



PROCESS(SYNTHESIZED_WIRE_68,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_69 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_69 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_68)) THEN
	SYNTHESIZED_WIRE_69 <= SYNTHESIZED_WIRE_34;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_34 <= NOT(SYNTHESIZED_WIRE_69);



PROCESS(SYNTHESIZED_WIRE_69,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_70 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_70 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_69)) THEN
	SYNTHESIZED_WIRE_70 <= SYNTHESIZED_WIRE_36;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_36 <= NOT(SYNTHESIZED_WIRE_70);



PROCESS(SYNTHESIZED_WIRE_70,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_71 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_71 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_70)) THEN
	SYNTHESIZED_WIRE_71 <= SYNTHESIZED_WIRE_38;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_38 <= NOT(SYNTHESIZED_WIRE_71);



PROCESS(SYNTHESIZED_WIRE_71,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_72 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_72 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_71)) THEN
	SYNTHESIZED_WIRE_72 <= SYNTHESIZED_WIRE_40;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_40 <= NOT(SYNTHESIZED_WIRE_72);



PROCESS(SYNTHESIZED_WIRE_72,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	clkOUT_ALTERA_SYNTHESIZED <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	clkOUT_ALTERA_SYNTHESIZED <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_72)) THEN
	clkOUT_ALTERA_SYNTHESIZED <= SYNTHESIZED_WIRE_42;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_67,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_73 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_73 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_67)) THEN
	SYNTHESIZED_WIRE_73 <= SYNTHESIZED_WIRE_44;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_42 <= NOT(clkOUT_ALTERA_SYNTHESIZED);



SYNTHESIZED_WIRE_44 <= NOT(SYNTHESIZED_WIRE_73);



PROCESS(SYNTHESIZED_WIRE_73,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_74 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_74 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_73)) THEN
	SYNTHESIZED_WIRE_74 <= SYNTHESIZED_WIRE_46;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_46 <= NOT(SYNTHESIZED_WIRE_74);



PROCESS(SYNTHESIZED_WIRE_74,rst,SYNTHESIZED_WIRE_50)
BEGIN
IF (rst = '0') THEN
	SYNTHESIZED_WIRE_52 <= '0';
ELSIF (SYNTHESIZED_WIRE_50 = '0') THEN
	SYNTHESIZED_WIRE_52 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_74)) THEN
	SYNTHESIZED_WIRE_52 <= SYNTHESIZED_WIRE_48;
END IF;
END PROCESS;

clkOUT <= clkOUT_ALTERA_SYNTHESIZED;

END bdf_type;